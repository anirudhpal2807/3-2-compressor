* File name: D:\cmos project\3_2_anirudhpal\3_2_anirudh.sch
* Software version: DSCH 2.7f
* Created 11/10/2024 11:43:33 PM
*
* Voltage and current sources
*
VBTN1 3 0 DC 0 PULSE(0 1.2 1.00N 0.1N 0.1N 1.00N 3.00N )
VBTN2 2 0 DC 0 PULSE(0 1.2 2.00N 0.1N 0.1N 2.00N 5.00N )
VBTN3 6 0 DC 0 PULSE(0 1.2 3.00N 0.1N 0.1N 3.00N 7.00N )
*
* Passive devices
*
*
* Active devices
*
MP1 1 2 10 1  W= L=
MP2 1 3 10 1  W= L=
MP3 1 10 5 1  W= L=
MN1 11 2 10 11  W= L=
MN2 0 3 11 0  W= L=
MN3 12 10 5 12  W= L=
MN4 0 2 12 0  W= L=
MN5 0 3 12 0  W= L=
MP4 1 2 13 1  W= L=
MP5 13 3 5 13  W= L=
MP6 1 5 4 1  W= L=
MN6 0 5 4 0  W= L=
MP7 1 6 14 1  W= L=
MP8 1 4 14 1  W= L=
MP9 1 14 8 1  W= L=
MN7 15 6 14 15  W= L=
MN8 0 4 15 0  W= L=
MN9 16 14 8 16  W= L=
MN10 0 6 16 0  W= L=
MN11 0 4 16 0  W= L=
MP10 1 6 17 1  W= L=
MP11 17 4 8 17  W= L=
MP12 1 8 7 1  W= L=
MN12 0 8 7 0  W= L=
*
* Warning: "spice.lib" not found, model not declared
.TRAN 0.1ns 250ns
*--Pspice--
.PROBE
.OPTIONS DELMIN=0 RELTOL=1E-6
.END
